// module subtract_32(x,y,out);
//     input [31:0] x;
//     input [31:0] y;
//     output [31:0] out;

//     not 0_bit(out[0], x[0], y[0]); 
//     not 1_bit(out[1], x[1], y[1]); 
//     not 2_bit(out[2], x[2], y[2]); 
//     not 3_bit(out[3], x[3], y[3]); 
//     not 4_bit(out[4], x[4], y[4]); 

//     not 5_bit(out[5], x[5], y[5]); 
//     not 6_bit(out[6], x[6], y[6]); 
//     not 7_bit(out[7], x[7], y[7]); 
//     not 8_bit(out[8], x[8], y[8]); 
//     not 9_bit(out[9], x[9], y[9]); 

//     not 10_bit(out[10], x[10], y[10]); 
//     not 11_bit(out[11], x[11], y[11]); 
//     not 12_bit(out[12], x[12], y[12]); 
//     not 13_bit(out[13], x[13], y[13]); 
//     not 14_bit(out[14], x[14], y[14]); 

//     not 15_bit(out[15], x[15], y[15]); 
//     not 16_bit(out[16], x[16], y[16]); 
//     not 17_bit(out[17], x[17], y[17]); 
//     not 18_bit(out[18], x[18], y[18]); 
//     not 19_bit(out[19], x[19], y[19]);

//     not 20_bit(out[20], x[20], y[20]); 
//     not 21_bit(out[21], x[21], y[21]); 
//     not 22_bit(out[22], x[22], y[22]); 
//     not 23_bit(out[23], x[23], y[23]); 
//     not 24_bit(out[24], x[24], y[24]);

//     not 25_bit(out[25], x[25], y[25]); 
//     not 26_bit(out[26], x[26], y[26]); 
//     not 27_bit(out[27], x[27], y[27]); 
//     not 28_bit(out[28], x[28], y[28]); 
//     not 29_bit(out[29], x[29], y[29]);

//     not 30_bit(out[30], x[30], y[30]); 
//     not 31_bit(out[31], x[31], y[31]);
    

// endmodule