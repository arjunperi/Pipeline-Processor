module not_32(x,out);
    input [31:0] x;
    output [31:0] out;

    not bit_0(out[0], x[0]); 
    not bit_1(out[1], x[1]); 
    not bit_2(out[2], x[2]); 
    not bit_3(out[3], x[3]); 
    not bit_4(out[4], x[4]); 

    not bit_5(out[5], x[5]); 
    not bit_6(out[6], x[6]); 
    not bit_7(out[7], x[7]); 
    not bit_8(out[8], x[8]); 
    not bit_9(out[9], x[9]); 

    not bit_10(out[10], x[10]); 
    not bit_11(out[11], x[11]); 
    not bit_12(out[12], x[12]); 
    not bit_13(out[13], x[13]); 
    not bit_14(out[14], x[14]); 

    not bit_15(out[15], x[15]); 
    not bit_16(out[16], x[16]); 
    not bit_17(out[17], x[17]); 
    not bit_18(out[18], x[18]); 
    not bit_19(out[19], x[19]);

    not bit_20(out[20], x[20]); 
    not bit_21(out[21], x[21]); 
    not bit_22(out[22], x[22]); 
    not bit_23(out[23], x[23]); 
    not bit_24(out[24], x[24]);

    not bit_25(out[25], x[25]); 
    not bit_26(out[26], x[26]); 
    not bit_27(out[27], x[27]); 
    not bit_28(out[28], x[28]); 
    not bit_29(out[29], x[29]);

    not bit_30(out[30], x[30]); 
    not bit_31(out[31], x[31]);
    

endmodule